module _ROM(Addr,Data);
	input [31:0] Addr;
	output [31:0] Data;
	
	reg [31:0] Data;

	always @(*)
		case(Addr[7:2])
			0: Data=32'b00001000010000000000000000000010;
			1: Data=32'b00001000010000000000000000001101;
			2: Data=32'b00111100000010010100000000000000;
			3: Data=32'b00111100000010100000000000010000;
			4: Data=32'b00000000000010100101010000000010;
			5: Data=32'b00000001001010100100100000100001;
			6: Data=32'b00111100000010100100000000000000;
			7: Data=32'b00111100000010110000000000001100;
			8: Data=32'b00000000000010110101110000000010;
			9: Data=32'b00000001010010110101000000100001;
			10: Data=32'b10001101001010110000000000000000;
			11: Data=32'b10101101010010110000000000000000;
			12: Data=32'b00001000010000000000000000000010;
			13: Data=32'b00001000010000000000000000000010;
		   default:	Data=32'h00000000;
		endcase
endmodule
